library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;
use IEEE.NUMERIC_STD.ALL;


PACKAGE parameter IS
  TYPE corrData IS ARRAY(0 TO 280) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
END PACKAGE;



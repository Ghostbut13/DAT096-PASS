
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.config_state_package.all;
use work.i2c_type_package.all;

entity Wrapper_ACFC_i2c_tb is
  
end entity Wrapper_ACFC_i2c_tb;

architecture arch of Wrapper_ACFC_i2c_tb is

  component Wrapper_ACFC_i2c is
    port (
      finish_config_input: in std_logic;
      -- config THE MODE
      I2S_mode          : in    std_logic;
      master_mode       : in    std_logic;
      GPIO_MCLK         : in    std_logic;
      FS_48k_256_BCLK   : in    std_logic;
      MCLK_root         : in    std_logic;

      -- MCLK(GPIO)-generated by PLL and SHDNZ
      SHDNZ             : out   std_logic;
      MCLK              : out   std_logic;

      -- clk and rstn
      clk               : in    std_logic;
      rstn              : in    std_logic;
      
      -- control ready
      SW_vdd_ok         : in    std_logic;
      SHDNZ_ready       : in    std_logic;
      
      -- FSYNC and BCLK 
      FSYNC             : out   std_logic;
      BCLK              : out   std_logic;
      
      -- i2c communication
      SDA               : inout std_logic;
      SCL               : out   std_logic
      
      );
  end component Wrapper_ACFC_i2c;

  signal clk_tb  : std_logic := '1';
  signal rstn_tb : std_logic := '1';
  signal SCL_tb  : std_logic;
  signal SDA_tb  : std_logic;
  signal SHDNZ_pin_tb : std_logic := '0';
  signal SW_vdd_ok_tb : std_logic := '0';
  signal finish_config_input_tb : std_logic := '0';



  ----------------------------------------
  signal FSYNC_tb :  std_logic ;

  signal I2S_mode_tb    :   std_logic := '0';
  signal master_mode_tb :   std_logic := '0';
  signal GPIO_MCLK_tb   :   std_logic := '0';
  signal FS_48k_256_BCLK_tb :std_logic := '0';
  signal MCLK_root_tb   :   std_logic := '0';
  ----------------------------------------
  
begin  -- architecture arch_I2C_master_for_temperature

  inst_W: Wrapper_ACFC_i2c
    port map (
      finish_config_input   => finish_config_input_tb,
      I2S_mode          => I2S_mode_tb,
      master_mode       => master_mode_tb,
      GPIO_MCLK         => GPIO_MCLK_tb  ,
      FS_48k_256_BCLK   => FS_48k_256_BCLK_tb,
      MCLK_root         => MCLK_root_tb,
      
      clk               => clk_tb,
      rstn              => rstn_tb,

      SW_vdd_ok         => SW_vdd_ok_tb,
      SHDNZ_ready       => SHDNZ_pin_tb,

      SDA => SDA_tb,
      SCL => SCL_tb,
      
      FSYNC             => FSYNC_tb
      );


  proc_clk_gen : 
  process
  begin
    wait for 5 ns;
    clk_tb <= not(clk_tb) ;
  end process proc_clk_gen;
  rstn_tb <= '0' after 1 ns,
             '1' after 2 ns;


  
  SW_vdd_ok_tb <= '1' after 243 ns;
                  -- '0' after when_can_done * 19 + 10 ns,
                  -- '1' after when_can_done * 22;

  SHDNZ_pin_tb <= '1' after 991 ns,
                  -- good 28 10 29
                  --'0' after when_can_done * 28 + 10 ns,
                  --'1' after when_can_done * 29;
                  -- fixed time : 14000000
                  '0' after (14000000 ns + 20000000 ns ),
                  '1' after (14600000 ns + 20000000 ns);

 
  ----------------------------------------
  -- I2S_mode_tb <= '1' after 10000000 ns,
  --                '0' after (300000 ns+10000000 ns);


  -- GPIO_MCLK_tb <= '1' after 11000000 ns,
  --                 '0' after (300000 ns+11000000 ns);

  -- master_mode_tb <= '1' after 12000000 ns,
  --                   '0' after (300000 ns+12000000 ns);

  -- FS_48k_256_BCLK_tb <= '1' after 13000000 ns,
  --                       '0' after (300000 ns+13000000 ns);
  ----------------------------------------


  finish_config_input_tb <= '1' after 16000000 ns;

  
  ----------------------------------------
  


  GPIO_MCLK_tb          <= '1' after 6000000 ns;
                           --'0' after 6000100 ns;

  master_mode_tb        <= '1' after 7300000 ns;
                           --'0' after 7300100 ns;
  
  FS_48k_256_BCLK_tb    <= '1' after 8300000 ns;
                           --'0' after 8300100 ns;
  
  I2S_mode_tb           <= '1' after 9300000 ns;
                           --'0' after 9300100 ns;
  
  MCLK_root_tb          <= '1' after 10300000 ns;
                           --'0' after 10301000 ns;
  
  
----------------------------------------
end architecture arch;

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

PACKAGE parameter IS
  CONSTANT SIGNAL_WIDTH :INTEGER := 16;
  CONSTANT REGISTER_LENGTH : INTEGER := 5;
  constant LEN_DATA: integer:=23;
  TYPE outputdata IS ARRAY(0 TO REGISTER_LENGTH-1) OF STD_LOGIC_VECTOR(SIGNAL_WIDTH-1 DOWNTO 0);
  TYPE testdata IS ARRAY(0 TO 4) OF STD_LOGIC_VECTOR(SIGNAL_WIDTH-1 DOWNTO 0);
  
  SIGNAL test_data: testdata :=("1010101010101010","0101010101010101","1111111100000000","0000000011111111","1111111111111111");
END PACKAGE;


-- ----------- -------------------------------------------------------------


LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE IEEE.numeric_std.ALL;

PACKAGE mlhdlc_aesd_fixpt_pkg IS
  TYPE vector_of_std_logic_vector8 IS ARRAY (NATURAL RANGE <>) OF std_logic_vector(7 DOWNTO 0);
  TYPE vector_of_unsigned8 IS ARRAY (NATURAL RANGE <>) OF unsigned(7 DOWNTO 0);
  TYPE vector_of_signed32 IS ARRAY (NATURAL RANGE <>) OF signed(31 DOWNTO 0);
  TYPE vector_of_signed16 IS ARRAY (NATURAL RANGE <>) OF signed(15 DOWNTO 0);
  TYPE vector_of_unsigned6 IS ARRAY (NATURAL RANGE <>) OF unsigned(5 DOWNTO 0);
  TYPE vector_of_unsigned5 IS ARRAY (NATURAL RANGE <>) OF unsigned(4 DOWNTO 0);
  TYPE vector_of_unsigned7 IS ARRAY (NATURAL RANGE <>) OF unsigned(6 DOWNTO 0);
  TYPE vector_of_unsigned9 IS ARRAY (NATURAL RANGE <>) OF unsigned(8 DOWNTO 0);
  

  CONSTANT cipherkey  : vector_of_unsigned8(0 TO 15) := (to_unsigned(16#6C#, 8), to_unsigned(16#EA#, 8), to_unsigned(16#CB#, 8), to_unsigned(16#F6#, 8), to_unsigned(16#A8#, 8), to_unsigned(16#09#, 8), to_unsigned(16#D9#, 8), to_unsigned(16#EF#, 8), to_unsigned(16#AE#, 8), to_unsigned(16#C2#, 8), to_unsigned(16#BE#, 8), to_unsigned(16#64#, 8), to_unsigned(16#A8#, 8), to_unsigned(16#2C#, 8), to_unsigned(16#B5#, 8), to_unsigned(16#08#,8));


 -- CONSTANT ciphertext  : vector_of_unsigned8(0 TO 15) := (to_unsigned(16#1F#, 8), to_unsigned(16#9D#, 8), to_unsigned(16#05#, 8), to_unsigned(16#17#, 8), to_unsigned(16#7B#, 8), to_unsigned(16#B0#, 8), to_unsigned(16#5F#, 8), to_unsigned(16#87#, 8), to_unsigned(16#99#, 8), to_unsigned(16#7A#, 8), to_unsigned(16#AE#, 8), to_unsigned(16#F3#, 8), to_unsigned(16#9E#, 8), to_unsigned(16#82#, 8), to_unsigned(16#51#, 8), to_unsigned(16#CC#,8));
 
  -- Constants
  CONSTANT tmp_3                          : vector_of_unsigned8(0 TO 255) := 
    (to_unsigned(16#63#, 8), to_unsigned(16#7C#, 8), to_unsigned(16#77#, 8), to_unsigned(16#7B#, 8),
     to_unsigned(16#F2#, 8), to_unsigned(16#6B#, 8), to_unsigned(16#6F#, 8), to_unsigned(16#C5#, 8),
     to_unsigned(16#30#, 8), to_unsigned(16#01#, 8), to_unsigned(16#67#, 8), to_unsigned(16#2B#, 8),
     to_unsigned(16#FE#, 8), to_unsigned(16#D7#, 8), to_unsigned(16#AB#, 8), to_unsigned(16#76#, 8),
     to_unsigned(16#CA#, 8), to_unsigned(16#82#, 8), to_unsigned(16#C9#, 8), to_unsigned(16#7D#, 8),
     to_unsigned(16#FA#, 8), to_unsigned(16#59#, 8), to_unsigned(16#47#, 8), to_unsigned(16#F0#, 8),
     to_unsigned(16#AD#, 8), to_unsigned(16#D4#, 8), to_unsigned(16#A2#, 8), to_unsigned(16#AF#, 8),
     to_unsigned(16#9C#, 8), to_unsigned(16#A4#, 8), to_unsigned(16#72#, 8), to_unsigned(16#C0#, 8),
     to_unsigned(16#B7#, 8), to_unsigned(16#FD#, 8), to_unsigned(16#93#, 8), to_unsigned(16#26#, 8),
     to_unsigned(16#36#, 8), to_unsigned(16#3F#, 8), to_unsigned(16#F7#, 8), to_unsigned(16#CC#, 8),
     to_unsigned(16#34#, 8), to_unsigned(16#A5#, 8), to_unsigned(16#E5#, 8), to_unsigned(16#F1#, 8),
     to_unsigned(16#71#, 8), to_unsigned(16#D8#, 8), to_unsigned(16#31#, 8), to_unsigned(16#15#, 8),
     to_unsigned(16#04#, 8), to_unsigned(16#C7#, 8), to_unsigned(16#23#, 8), to_unsigned(16#C3#, 8),
     to_unsigned(16#18#, 8), to_unsigned(16#96#, 8), to_unsigned(16#05#, 8), to_unsigned(16#9A#, 8),
     to_unsigned(16#07#, 8), to_unsigned(16#12#, 8), to_unsigned(16#80#, 8), to_unsigned(16#E2#, 8),
     to_unsigned(16#EB#, 8), to_unsigned(16#27#, 8), to_unsigned(16#B2#, 8), to_unsigned(16#75#, 8),
     to_unsigned(16#09#, 8), to_unsigned(16#83#, 8), to_unsigned(16#2C#, 8), to_unsigned(16#1A#, 8),
     to_unsigned(16#1B#, 8), to_unsigned(16#6E#, 8), to_unsigned(16#5A#, 8), to_unsigned(16#A0#, 8),
     to_unsigned(16#52#, 8), to_unsigned(16#3B#, 8), to_unsigned(16#D6#, 8), to_unsigned(16#B3#, 8),
     to_unsigned(16#29#, 8), to_unsigned(16#E3#, 8), to_unsigned(16#2F#, 8), to_unsigned(16#84#, 8),
     to_unsigned(16#53#, 8), to_unsigned(16#D1#, 8), to_unsigned(16#00#, 8), to_unsigned(16#ED#, 8),
     to_unsigned(16#20#, 8), to_unsigned(16#FC#, 8), to_unsigned(16#B1#, 8), to_unsigned(16#5B#, 8),
     to_unsigned(16#6A#, 8), to_unsigned(16#CB#, 8), to_unsigned(16#BE#, 8), to_unsigned(16#39#, 8),
     to_unsigned(16#4A#, 8), to_unsigned(16#4C#, 8), to_unsigned(16#58#, 8), to_unsigned(16#CF#, 8),
     to_unsigned(16#D0#, 8), to_unsigned(16#EF#, 8), to_unsigned(16#AA#, 8), to_unsigned(16#FB#, 8),
     to_unsigned(16#43#, 8), to_unsigned(16#4D#, 8), to_unsigned(16#33#, 8), to_unsigned(16#85#, 8),
     to_unsigned(16#45#, 8), to_unsigned(16#F9#, 8), to_unsigned(16#02#, 8), to_unsigned(16#7F#, 8),
     to_unsigned(16#50#, 8), to_unsigned(16#3C#, 8), to_unsigned(16#9F#, 8), to_unsigned(16#A8#, 8),
     to_unsigned(16#51#, 8), to_unsigned(16#A3#, 8), to_unsigned(16#40#, 8), to_unsigned(16#8F#, 8),
     to_unsigned(16#92#, 8), to_unsigned(16#9D#, 8), to_unsigned(16#38#, 8), to_unsigned(16#F5#, 8),
     to_unsigned(16#BC#, 8), to_unsigned(16#B6#, 8), to_unsigned(16#DA#, 8), to_unsigned(16#21#, 8),
     to_unsigned(16#10#, 8), to_unsigned(16#FF#, 8), to_unsigned(16#F3#, 8), to_unsigned(16#D2#, 8),
     to_unsigned(16#CD#, 8), to_unsigned(16#0C#, 8), to_unsigned(16#13#, 8), to_unsigned(16#EC#, 8),
     to_unsigned(16#5F#, 8), to_unsigned(16#97#, 8), to_unsigned(16#44#, 8), to_unsigned(16#17#, 8),
     to_unsigned(16#C4#, 8), to_unsigned(16#A7#, 8), to_unsigned(16#7E#, 8), to_unsigned(16#3D#, 8),
     to_unsigned(16#64#, 8), to_unsigned(16#5D#, 8), to_unsigned(16#19#, 8), to_unsigned(16#73#, 8),
     to_unsigned(16#60#, 8), to_unsigned(16#81#, 8), to_unsigned(16#4F#, 8), to_unsigned(16#DC#, 8),
     to_unsigned(16#22#, 8), to_unsigned(16#2A#, 8), to_unsigned(16#90#, 8), to_unsigned(16#88#, 8),
     to_unsigned(16#46#, 8), to_unsigned(16#EE#, 8), to_unsigned(16#B8#, 8), to_unsigned(16#14#, 8),
     to_unsigned(16#DE#, 8), to_unsigned(16#5E#, 8), to_unsigned(16#0B#, 8), to_unsigned(16#DB#, 8),
     to_unsigned(16#E0#, 8), to_unsigned(16#32#, 8), to_unsigned(16#3A#, 8), to_unsigned(16#0A#, 8),
     to_unsigned(16#49#, 8), to_unsigned(16#06#, 8), to_unsigned(16#24#, 8), to_unsigned(16#5C#, 8),
     to_unsigned(16#C2#, 8), to_unsigned(16#D3#, 8), to_unsigned(16#AC#, 8), to_unsigned(16#62#, 8),
     to_unsigned(16#91#, 8), to_unsigned(16#95#, 8), to_unsigned(16#E4#, 8), to_unsigned(16#79#, 8),
     to_unsigned(16#E7#, 8), to_unsigned(16#C8#, 8), to_unsigned(16#37#, 8), to_unsigned(16#6D#, 8),
     to_unsigned(16#8D#, 8), to_unsigned(16#D5#, 8), to_unsigned(16#4E#, 8), to_unsigned(16#A9#, 8),
     to_unsigned(16#6C#, 8), to_unsigned(16#56#, 8), to_unsigned(16#F4#, 8), to_unsigned(16#EA#, 8),
     to_unsigned(16#65#, 8), to_unsigned(16#7A#, 8), to_unsigned(16#AE#, 8), to_unsigned(16#08#, 8),
     to_unsigned(16#BA#, 8), to_unsigned(16#78#, 8), to_unsigned(16#25#, 8), to_unsigned(16#2E#, 8),
     to_unsigned(16#1C#, 8), to_unsigned(16#A6#, 8), to_unsigned(16#B4#, 8), to_unsigned(16#C6#, 8),
     to_unsigned(16#E8#, 8), to_unsigned(16#DD#, 8), to_unsigned(16#74#, 8), to_unsigned(16#1F#, 8),
     to_unsigned(16#4B#, 8), to_unsigned(16#BD#, 8), to_unsigned(16#8B#, 8), to_unsigned(16#8A#, 8),
     to_unsigned(16#70#, 8), to_unsigned(16#3E#, 8), to_unsigned(16#B5#, 8), to_unsigned(16#66#, 8),
     to_unsigned(16#48#, 8), to_unsigned(16#03#, 8), to_unsigned(16#F6#, 8), to_unsigned(16#0E#, 8),
     to_unsigned(16#61#, 8), to_unsigned(16#35#, 8), to_unsigned(16#57#, 8), to_unsigned(16#B9#, 8),
     to_unsigned(16#86#, 8), to_unsigned(16#C1#, 8), to_unsigned(16#1D#, 8), to_unsigned(16#9E#, 8),
     to_unsigned(16#E1#, 8), to_unsigned(16#F8#, 8), to_unsigned(16#98#, 8), to_unsigned(16#11#, 8),
     to_unsigned(16#69#, 8), to_unsigned(16#D9#, 8), to_unsigned(16#8E#, 8), to_unsigned(16#94#, 8),
     to_unsigned(16#9B#, 8), to_unsigned(16#1E#, 8), to_unsigned(16#87#, 8), to_unsigned(16#E9#, 8),
     to_unsigned(16#CE#, 8), to_unsigned(16#55#, 8), to_unsigned(16#28#, 8), to_unsigned(16#DF#, 8),
     to_unsigned(16#8C#, 8), to_unsigned(16#A1#, 8), to_unsigned(16#89#, 8), to_unsigned(16#0D#, 8),
     to_unsigned(16#BF#, 8), to_unsigned(16#E6#, 8), to_unsigned(16#42#, 8), to_unsigned(16#68#, 8),
     to_unsigned(16#41#, 8), to_unsigned(16#99#, 8), to_unsigned(16#2D#, 8), to_unsigned(16#0F#, 8),
     to_unsigned(16#B0#, 8), to_unsigned(16#54#, 8), to_unsigned(16#BB#, 8), to_unsigned(16#16#, 8));  -- ufix8 [256]
  CONSTANT nc                             : vector_of_unsigned8(0 TO 255) := 
    (to_unsigned(16#63#, 8), to_unsigned(16#7C#, 8), to_unsigned(16#77#, 8), to_unsigned(16#7B#, 8),
     to_unsigned(16#F2#, 8), to_unsigned(16#6B#, 8), to_unsigned(16#6F#, 8), to_unsigned(16#C5#, 8),
     to_unsigned(16#30#, 8), to_unsigned(16#01#, 8), to_unsigned(16#67#, 8), to_unsigned(16#2B#, 8),
     to_unsigned(16#FE#, 8), to_unsigned(16#D7#, 8), to_unsigned(16#AB#, 8), to_unsigned(16#76#, 8),
     to_unsigned(16#CA#, 8), to_unsigned(16#82#, 8), to_unsigned(16#C9#, 8), to_unsigned(16#7D#, 8),
     to_unsigned(16#FA#, 8), to_unsigned(16#59#, 8), to_unsigned(16#47#, 8), to_unsigned(16#F0#, 8),
     to_unsigned(16#AD#, 8), to_unsigned(16#D4#, 8), to_unsigned(16#A2#, 8), to_unsigned(16#AF#, 8),
     to_unsigned(16#9C#, 8), to_unsigned(16#A4#, 8), to_unsigned(16#72#, 8), to_unsigned(16#C0#, 8),
     to_unsigned(16#B7#, 8), to_unsigned(16#FD#, 8), to_unsigned(16#93#, 8), to_unsigned(16#26#, 8),
     to_unsigned(16#36#, 8), to_unsigned(16#3F#, 8), to_unsigned(16#F7#, 8), to_unsigned(16#CC#, 8),
     to_unsigned(16#34#, 8), to_unsigned(16#A5#, 8), to_unsigned(16#E5#, 8), to_unsigned(16#F1#, 8),
     to_unsigned(16#71#, 8), to_unsigned(16#D8#, 8), to_unsigned(16#31#, 8), to_unsigned(16#15#, 8),
     to_unsigned(16#04#, 8), to_unsigned(16#C7#, 8), to_unsigned(16#23#, 8), to_unsigned(16#C3#, 8),
     to_unsigned(16#18#, 8), to_unsigned(16#96#, 8), to_unsigned(16#05#, 8), to_unsigned(16#9A#, 8),
     to_unsigned(16#07#, 8), to_unsigned(16#12#, 8), to_unsigned(16#80#, 8), to_unsigned(16#E2#, 8),
     to_unsigned(16#EB#, 8), to_unsigned(16#27#, 8), to_unsigned(16#B2#, 8), to_unsigned(16#75#, 8),
     to_unsigned(16#09#, 8), to_unsigned(16#83#, 8), to_unsigned(16#2C#, 8), to_unsigned(16#1A#, 8),
     to_unsigned(16#1B#, 8), to_unsigned(16#6E#, 8), to_unsigned(16#5A#, 8), to_unsigned(16#A0#, 8),
     to_unsigned(16#52#, 8), to_unsigned(16#3B#, 8), to_unsigned(16#D6#, 8), to_unsigned(16#B3#, 8),
     to_unsigned(16#29#, 8), to_unsigned(16#E3#, 8), to_unsigned(16#2F#, 8), to_unsigned(16#84#, 8),
     to_unsigned(16#53#, 8), to_unsigned(16#D1#, 8), to_unsigned(16#00#, 8), to_unsigned(16#ED#, 8),
     to_unsigned(16#20#, 8), to_unsigned(16#FC#, 8), to_unsigned(16#B1#, 8), to_unsigned(16#5B#, 8),
     to_unsigned(16#6A#, 8), to_unsigned(16#CB#, 8), to_unsigned(16#BE#, 8), to_unsigned(16#39#, 8),
     to_unsigned(16#4A#, 8), to_unsigned(16#4C#, 8), to_unsigned(16#58#, 8), to_unsigned(16#CF#, 8),
     to_unsigned(16#D0#, 8), to_unsigned(16#EF#, 8), to_unsigned(16#AA#, 8), to_unsigned(16#FB#, 8),
     to_unsigned(16#43#, 8), to_unsigned(16#4D#, 8), to_unsigned(16#33#, 8), to_unsigned(16#85#, 8),
     to_unsigned(16#45#, 8), to_unsigned(16#F9#, 8), to_unsigned(16#02#, 8), to_unsigned(16#7F#, 8),
     to_unsigned(16#50#, 8), to_unsigned(16#3C#, 8), to_unsigned(16#9F#, 8), to_unsigned(16#A8#, 8),
     to_unsigned(16#51#, 8), to_unsigned(16#A3#, 8), to_unsigned(16#40#, 8), to_unsigned(16#8F#, 8),
     to_unsigned(16#92#, 8), to_unsigned(16#9D#, 8), to_unsigned(16#38#, 8), to_unsigned(16#F5#, 8),
     to_unsigned(16#BC#, 8), to_unsigned(16#B6#, 8), to_unsigned(16#DA#, 8), to_unsigned(16#21#, 8),
     to_unsigned(16#10#, 8), to_unsigned(16#FF#, 8), to_unsigned(16#F3#, 8), to_unsigned(16#D2#, 8),
     to_unsigned(16#CD#, 8), to_unsigned(16#0C#, 8), to_unsigned(16#13#, 8), to_unsigned(16#EC#, 8),
     to_unsigned(16#5F#, 8), to_unsigned(16#97#, 8), to_unsigned(16#44#, 8), to_unsigned(16#17#, 8),
     to_unsigned(16#C4#, 8), to_unsigned(16#A7#, 8), to_unsigned(16#7E#, 8), to_unsigned(16#3D#, 8),
     to_unsigned(16#64#, 8), to_unsigned(16#5D#, 8), to_unsigned(16#19#, 8), to_unsigned(16#73#, 8),
     to_unsigned(16#60#, 8), to_unsigned(16#81#, 8), to_unsigned(16#4F#, 8), to_unsigned(16#DC#, 8),
     to_unsigned(16#22#, 8), to_unsigned(16#2A#, 8), to_unsigned(16#90#, 8), to_unsigned(16#88#, 8),
     to_unsigned(16#46#, 8), to_unsigned(16#EE#, 8), to_unsigned(16#B8#, 8), to_unsigned(16#14#, 8),
     to_unsigned(16#DE#, 8), to_unsigned(16#5E#, 8), to_unsigned(16#0B#, 8), to_unsigned(16#DB#, 8),
     to_unsigned(16#E0#, 8), to_unsigned(16#32#, 8), to_unsigned(16#3A#, 8), to_unsigned(16#0A#, 8),
     to_unsigned(16#49#, 8), to_unsigned(16#06#, 8), to_unsigned(16#24#, 8), to_unsigned(16#5C#, 8),
     to_unsigned(16#C2#, 8), to_unsigned(16#D3#, 8), to_unsigned(16#AC#, 8), to_unsigned(16#62#, 8),
     to_unsigned(16#91#, 8), to_unsigned(16#95#, 8), to_unsigned(16#E4#, 8), to_unsigned(16#79#, 8),
     to_unsigned(16#E7#, 8), to_unsigned(16#C8#, 8), to_unsigned(16#37#, 8), to_unsigned(16#6D#, 8),
     to_unsigned(16#8D#, 8), to_unsigned(16#D5#, 8), to_unsigned(16#4E#, 8), to_unsigned(16#A9#, 8),
     to_unsigned(16#6C#, 8), to_unsigned(16#56#, 8), to_unsigned(16#F4#, 8), to_unsigned(16#EA#, 8),
     to_unsigned(16#65#, 8), to_unsigned(16#7A#, 8), to_unsigned(16#AE#, 8), to_unsigned(16#08#, 8),
     to_unsigned(16#BA#, 8), to_unsigned(16#78#, 8), to_unsigned(16#25#, 8), to_unsigned(16#2E#, 8),
     to_unsigned(16#1C#, 8), to_unsigned(16#A6#, 8), to_unsigned(16#B4#, 8), to_unsigned(16#C6#, 8),
     to_unsigned(16#E8#, 8), to_unsigned(16#DD#, 8), to_unsigned(16#74#, 8), to_unsigned(16#1F#, 8),
     to_unsigned(16#4B#, 8), to_unsigned(16#BD#, 8), to_unsigned(16#8B#, 8), to_unsigned(16#8A#, 8),
     to_unsigned(16#70#, 8), to_unsigned(16#3E#, 8), to_unsigned(16#B5#, 8), to_unsigned(16#66#, 8),
     to_unsigned(16#48#, 8), to_unsigned(16#03#, 8), to_unsigned(16#F6#, 8), to_unsigned(16#0E#, 8),
     to_unsigned(16#61#, 8), to_unsigned(16#35#, 8), to_unsigned(16#57#, 8), to_unsigned(16#B9#, 8),
     to_unsigned(16#86#, 8), to_unsigned(16#C1#, 8), to_unsigned(16#1D#, 8), to_unsigned(16#9E#, 8),
     to_unsigned(16#E1#, 8), to_unsigned(16#F8#, 8), to_unsigned(16#98#, 8), to_unsigned(16#11#, 8),
     to_unsigned(16#69#, 8), to_unsigned(16#D9#, 8), to_unsigned(16#8E#, 8), to_unsigned(16#94#, 8),
     to_unsigned(16#9B#, 8), to_unsigned(16#1E#, 8), to_unsigned(16#87#, 8), to_unsigned(16#E9#, 8),
     to_unsigned(16#CE#, 8), to_unsigned(16#55#, 8), to_unsigned(16#28#, 8), to_unsigned(16#DF#, 8),
     to_unsigned(16#8C#, 8), to_unsigned(16#A1#, 8), to_unsigned(16#89#, 8), to_unsigned(16#0D#, 8),
     to_unsigned(16#BF#, 8), to_unsigned(16#E6#, 8), to_unsigned(16#42#, 8), to_unsigned(16#68#, 8),
     to_unsigned(16#41#, 8), to_unsigned(16#99#, 8), to_unsigned(16#2D#, 8), to_unsigned(16#0F#, 8),
     to_unsigned(16#B0#, 8), to_unsigned(16#54#, 8), to_unsigned(16#BB#, 8), to_unsigned(16#16#, 8));  -- ufix8 [256]
  CONSTANT nc_0                           : vector_of_unsigned8(0 TO 254) := 
    (to_unsigned(16#8D#, 8), to_unsigned(16#01#, 8), to_unsigned(16#02#, 8), to_unsigned(16#04#, 8),
     to_unsigned(16#08#, 8), to_unsigned(16#10#, 8), to_unsigned(16#20#, 8), to_unsigned(16#40#, 8),
     to_unsigned(16#80#, 8), to_unsigned(16#1B#, 8), to_unsigned(16#36#, 8), to_unsigned(16#6C#, 8),
     to_unsigned(16#D8#, 8), to_unsigned(16#AB#, 8), to_unsigned(16#4D#, 8), to_unsigned(16#9A#, 8),
     to_unsigned(16#2F#, 8), to_unsigned(16#5E#, 8), to_unsigned(16#BC#, 8), to_unsigned(16#63#, 8),
     to_unsigned(16#C6#, 8), to_unsigned(16#97#, 8), to_unsigned(16#35#, 8), to_unsigned(16#6A#, 8),
     to_unsigned(16#D4#, 8), to_unsigned(16#B3#, 8), to_unsigned(16#7D#, 8), to_unsigned(16#FA#, 8),
     to_unsigned(16#EF#, 8), to_unsigned(16#C5#, 8), to_unsigned(16#91#, 8), to_unsigned(16#39#, 8),
     to_unsigned(16#72#, 8), to_unsigned(16#E4#, 8), to_unsigned(16#D3#, 8), to_unsigned(16#BD#, 8),
     to_unsigned(16#61#, 8), to_unsigned(16#C2#, 8), to_unsigned(16#9F#, 8), to_unsigned(16#25#, 8),
     to_unsigned(16#4A#, 8), to_unsigned(16#94#, 8), to_unsigned(16#33#, 8), to_unsigned(16#66#, 8),
     to_unsigned(16#CC#, 8), to_unsigned(16#83#, 8), to_unsigned(16#1D#, 8), to_unsigned(16#3A#, 8),
     to_unsigned(16#74#, 8), to_unsigned(16#E8#, 8), to_unsigned(16#CB#, 8), to_unsigned(16#8D#, 8),
     to_unsigned(16#01#, 8), to_unsigned(16#02#, 8), to_unsigned(16#04#, 8), to_unsigned(16#08#, 8),
     to_unsigned(16#10#, 8), to_unsigned(16#20#, 8), to_unsigned(16#40#, 8), to_unsigned(16#80#, 8),
     to_unsigned(16#1B#, 8), to_unsigned(16#36#, 8), to_unsigned(16#6C#, 8), to_unsigned(16#D8#, 8),
     to_unsigned(16#AB#, 8), to_unsigned(16#4D#, 8), to_unsigned(16#9A#, 8), to_unsigned(16#2F#, 8),
     to_unsigned(16#5E#, 8), to_unsigned(16#BC#, 8), to_unsigned(16#63#, 8), to_unsigned(16#C6#, 8),
     to_unsigned(16#97#, 8), to_unsigned(16#35#, 8), to_unsigned(16#6A#, 8), to_unsigned(16#D4#, 8),
     to_unsigned(16#B3#, 8), to_unsigned(16#7D#, 8), to_unsigned(16#FA#, 8), to_unsigned(16#EF#, 8),
     to_unsigned(16#C5#, 8), to_unsigned(16#91#, 8), to_unsigned(16#39#, 8), to_unsigned(16#72#, 8),
     to_unsigned(16#E4#, 8), to_unsigned(16#D3#, 8), to_unsigned(16#BD#, 8), to_unsigned(16#61#, 8),
     to_unsigned(16#C2#, 8), to_unsigned(16#9F#, 8), to_unsigned(16#25#, 8), to_unsigned(16#4A#, 8),
     to_unsigned(16#94#, 8), to_unsigned(16#33#, 8), to_unsigned(16#66#, 8), to_unsigned(16#CC#, 8),
     to_unsigned(16#83#, 8), to_unsigned(16#1D#, 8), to_unsigned(16#3A#, 8), to_unsigned(16#74#, 8),
     to_unsigned(16#E8#, 8), to_unsigned(16#CB#, 8), to_unsigned(16#8D#, 8), to_unsigned(16#01#, 8),
     to_unsigned(16#02#, 8), to_unsigned(16#04#, 8), to_unsigned(16#08#, 8), to_unsigned(16#10#, 8),
     to_unsigned(16#20#, 8), to_unsigned(16#40#, 8), to_unsigned(16#80#, 8), to_unsigned(16#1B#, 8),
     to_unsigned(16#36#, 8), to_unsigned(16#6C#, 8), to_unsigned(16#D8#, 8), to_unsigned(16#AB#, 8),
     to_unsigned(16#4D#, 8), to_unsigned(16#9A#, 8), to_unsigned(16#2F#, 8), to_unsigned(16#5E#, 8),
     to_unsigned(16#BC#, 8), to_unsigned(16#63#, 8), to_unsigned(16#C6#, 8), to_unsigned(16#97#, 8),
     to_unsigned(16#35#, 8), to_unsigned(16#6A#, 8), to_unsigned(16#D4#, 8), to_unsigned(16#B3#, 8),
     to_unsigned(16#7D#, 8), to_unsigned(16#FA#, 8), to_unsigned(16#EF#, 8), to_unsigned(16#C5#, 8),
     to_unsigned(16#91#, 8), to_unsigned(16#39#, 8), to_unsigned(16#72#, 8), to_unsigned(16#E4#, 8),
     to_unsigned(16#D3#, 8), to_unsigned(16#BD#, 8), to_unsigned(16#61#, 8), to_unsigned(16#C2#, 8),
     to_unsigned(16#9F#, 8), to_unsigned(16#25#, 8), to_unsigned(16#4A#, 8), to_unsigned(16#94#, 8),
     to_unsigned(16#33#, 8), to_unsigned(16#66#, 8), to_unsigned(16#CC#, 8), to_unsigned(16#83#, 8),
     to_unsigned(16#1D#, 8), to_unsigned(16#3A#, 8), to_unsigned(16#74#, 8), to_unsigned(16#E8#, 8),
     to_unsigned(16#CB#, 8), to_unsigned(16#8D#, 8), to_unsigned(16#01#, 8), to_unsigned(16#02#, 8),
     to_unsigned(16#04#, 8), to_unsigned(16#08#, 8), to_unsigned(16#10#, 8), to_unsigned(16#20#, 8),
     to_unsigned(16#40#, 8), to_unsigned(16#80#, 8), to_unsigned(16#1B#, 8), to_unsigned(16#36#, 8),
     to_unsigned(16#6C#, 8), to_unsigned(16#D8#, 8), to_unsigned(16#AB#, 8), to_unsigned(16#4D#, 8),
     to_unsigned(16#9A#, 8), to_unsigned(16#2F#, 8), to_unsigned(16#5E#, 8), to_unsigned(16#BC#, 8),
     to_unsigned(16#63#, 8), to_unsigned(16#C6#, 8), to_unsigned(16#97#, 8), to_unsigned(16#35#, 8),
     to_unsigned(16#6A#, 8), to_unsigned(16#D4#, 8), to_unsigned(16#B3#, 8), to_unsigned(16#7D#, 8),
     to_unsigned(16#FA#, 8), to_unsigned(16#EF#, 8), to_unsigned(16#C5#, 8), to_unsigned(16#91#, 8),
     to_unsigned(16#39#, 8), to_unsigned(16#72#, 8), to_unsigned(16#E4#, 8), to_unsigned(16#D3#, 8),
     to_unsigned(16#BD#, 8), to_unsigned(16#61#, 8), to_unsigned(16#C2#, 8), to_unsigned(16#9F#, 8),
     to_unsigned(16#25#, 8), to_unsigned(16#4A#, 8), to_unsigned(16#94#, 8), to_unsigned(16#33#, 8),
     to_unsigned(16#66#, 8), to_unsigned(16#CC#, 8), to_unsigned(16#83#, 8), to_unsigned(16#1D#, 8),
     to_unsigned(16#3A#, 8), to_unsigned(16#74#, 8), to_unsigned(16#E8#, 8), to_unsigned(16#CB#, 8),
     to_unsigned(16#8D#, 8), to_unsigned(16#01#, 8), to_unsigned(16#02#, 8), to_unsigned(16#04#, 8),
     to_unsigned(16#08#, 8), to_unsigned(16#10#, 8), to_unsigned(16#20#, 8), to_unsigned(16#40#, 8),
     to_unsigned(16#80#, 8), to_unsigned(16#1B#, 8), to_unsigned(16#36#, 8), to_unsigned(16#6C#, 8),
     to_unsigned(16#D8#, 8), to_unsigned(16#AB#, 8), to_unsigned(16#4D#, 8), to_unsigned(16#9A#, 8),
     to_unsigned(16#2F#, 8), to_unsigned(16#5E#, 8), to_unsigned(16#BC#, 8), to_unsigned(16#63#, 8),
     to_unsigned(16#C6#, 8), to_unsigned(16#97#, 8), to_unsigned(16#35#, 8), to_unsigned(16#6A#, 8),
     to_unsigned(16#D4#, 8), to_unsigned(16#B3#, 8), to_unsigned(16#7D#, 8), to_unsigned(16#FA#, 8),
     to_unsigned(16#EF#, 8), to_unsigned(16#C5#, 8), to_unsigned(16#91#, 8), to_unsigned(16#39#, 8),
     to_unsigned(16#72#, 8), to_unsigned(16#E4#, 8), to_unsigned(16#D3#, 8), to_unsigned(16#BD#, 8),
     to_unsigned(16#61#, 8), to_unsigned(16#C2#, 8), to_unsigned(16#9F#, 8), to_unsigned(16#25#, 8),
     to_unsigned(16#4A#, 8), to_unsigned(16#94#, 8), to_unsigned(16#33#, 8), to_unsigned(16#66#, 8),
     to_unsigned(16#CC#, 8), to_unsigned(16#83#, 8), to_unsigned(16#1D#, 8), to_unsigned(16#3A#, 8),
     to_unsigned(16#74#, 8), to_unsigned(16#E8#, 8), to_unsigned(16#CB#, 8));  -- ufix8 [255]
  CONSTANT nc_2                           : vector_of_unsigned8(0 TO 255) := 
    (to_unsigned(16#52#, 8), to_unsigned(16#09#, 8), to_unsigned(16#6A#, 8), to_unsigned(16#D5#, 8),
     to_unsigned(16#30#, 8), to_unsigned(16#36#, 8), to_unsigned(16#A5#, 8), to_unsigned(16#38#, 8),
     to_unsigned(16#BF#, 8), to_unsigned(16#40#, 8), to_unsigned(16#A3#, 8), to_unsigned(16#9E#, 8),
     to_unsigned(16#81#, 8), to_unsigned(16#F3#, 8), to_unsigned(16#D7#, 8), to_unsigned(16#FB#, 8),
     to_unsigned(16#7C#, 8), to_unsigned(16#E3#, 8), to_unsigned(16#39#, 8), to_unsigned(16#82#, 8),
     to_unsigned(16#9B#, 8), to_unsigned(16#2F#, 8), to_unsigned(16#FF#, 8), to_unsigned(16#87#, 8),
     to_unsigned(16#34#, 8), to_unsigned(16#8E#, 8), to_unsigned(16#43#, 8), to_unsigned(16#44#, 8),
     to_unsigned(16#C4#, 8), to_unsigned(16#DE#, 8), to_unsigned(16#E9#, 8), to_unsigned(16#CB#, 8),
     to_unsigned(16#54#, 8), to_unsigned(16#7B#, 8), to_unsigned(16#94#, 8), to_unsigned(16#32#, 8),
     to_unsigned(16#A6#, 8), to_unsigned(16#C2#, 8), to_unsigned(16#23#, 8), to_unsigned(16#3D#, 8),
     to_unsigned(16#EE#, 8), to_unsigned(16#4C#, 8), to_unsigned(16#95#, 8), to_unsigned(16#0B#, 8),
     to_unsigned(16#42#, 8), to_unsigned(16#FA#, 8), to_unsigned(16#C3#, 8), to_unsigned(16#4E#, 8),
     to_unsigned(16#08#, 8), to_unsigned(16#2E#, 8), to_unsigned(16#A1#, 8), to_unsigned(16#66#, 8),
     to_unsigned(16#28#, 8), to_unsigned(16#D9#, 8), to_unsigned(16#24#, 8), to_unsigned(16#B2#, 8),
     to_unsigned(16#76#, 8), to_unsigned(16#5B#, 8), to_unsigned(16#A2#, 8), to_unsigned(16#49#, 8),
     to_unsigned(16#6D#, 8), to_unsigned(16#8B#, 8), to_unsigned(16#D1#, 8), to_unsigned(16#25#, 8),
     to_unsigned(16#72#, 8), to_unsigned(16#F8#, 8), to_unsigned(16#F6#, 8), to_unsigned(16#64#, 8),
     to_unsigned(16#86#, 8), to_unsigned(16#68#, 8), to_unsigned(16#98#, 8), to_unsigned(16#16#, 8),
     to_unsigned(16#D4#, 8), to_unsigned(16#A4#, 8), to_unsigned(16#5C#, 8), to_unsigned(16#CC#, 8),
     to_unsigned(16#5D#, 8), to_unsigned(16#65#, 8), to_unsigned(16#B6#, 8), to_unsigned(16#92#, 8),
     to_unsigned(16#6C#, 8), to_unsigned(16#70#, 8), to_unsigned(16#48#, 8), to_unsigned(16#50#, 8),
     to_unsigned(16#FD#, 8), to_unsigned(16#ED#, 8), to_unsigned(16#B9#, 8), to_unsigned(16#DA#, 8),
     to_unsigned(16#5E#, 8), to_unsigned(16#15#, 8), to_unsigned(16#46#, 8), to_unsigned(16#57#, 8),
     to_unsigned(16#A7#, 8), to_unsigned(16#8D#, 8), to_unsigned(16#9D#, 8), to_unsigned(16#84#, 8),
     to_unsigned(16#90#, 8), to_unsigned(16#D8#, 8), to_unsigned(16#AB#, 8), to_unsigned(16#00#, 8),
     to_unsigned(16#8C#, 8), to_unsigned(16#BC#, 8), to_unsigned(16#D3#, 8), to_unsigned(16#0A#, 8),
     to_unsigned(16#F7#, 8), to_unsigned(16#E4#, 8), to_unsigned(16#58#, 8), to_unsigned(16#05#, 8),
     to_unsigned(16#B8#, 8), to_unsigned(16#B3#, 8), to_unsigned(16#45#, 8), to_unsigned(16#06#, 8),
     to_unsigned(16#D0#, 8), to_unsigned(16#2C#, 8), to_unsigned(16#1E#, 8), to_unsigned(16#8F#, 8),
     to_unsigned(16#CA#, 8), to_unsigned(16#3F#, 8), to_unsigned(16#0F#, 8), to_unsigned(16#02#, 8),
     to_unsigned(16#C1#, 8), to_unsigned(16#AF#, 8), to_unsigned(16#BD#, 8), to_unsigned(16#03#, 8),
     to_unsigned(16#01#, 8), to_unsigned(16#13#, 8), to_unsigned(16#8A#, 8), to_unsigned(16#6B#, 8),
     to_unsigned(16#3A#, 8), to_unsigned(16#91#, 8), to_unsigned(16#11#, 8), to_unsigned(16#41#, 8),
     to_unsigned(16#4F#, 8), to_unsigned(16#67#, 8), to_unsigned(16#DC#, 8), to_unsigned(16#EA#, 8),
     to_unsigned(16#97#, 8), to_unsigned(16#F2#, 8), to_unsigned(16#CF#, 8), to_unsigned(16#CE#, 8),
     to_unsigned(16#F0#, 8), to_unsigned(16#B4#, 8), to_unsigned(16#E6#, 8), to_unsigned(16#73#, 8),
     to_unsigned(16#96#, 8), to_unsigned(16#AC#, 8), to_unsigned(16#74#, 8), to_unsigned(16#22#, 8),
     to_unsigned(16#E7#, 8), to_unsigned(16#AD#, 8), to_unsigned(16#35#, 8), to_unsigned(16#85#, 8),
     to_unsigned(16#E2#, 8), to_unsigned(16#F9#, 8), to_unsigned(16#37#, 8), to_unsigned(16#E8#, 8),
     to_unsigned(16#1C#, 8), to_unsigned(16#75#, 8), to_unsigned(16#DF#, 8), to_unsigned(16#6E#, 8),
     to_unsigned(16#47#, 8), to_unsigned(16#F1#, 8), to_unsigned(16#1A#, 8), to_unsigned(16#71#, 8),
     to_unsigned(16#1D#, 8), to_unsigned(16#29#, 8), to_unsigned(16#C5#, 8), to_unsigned(16#89#, 8),
     to_unsigned(16#6F#, 8), to_unsigned(16#B7#, 8), to_unsigned(16#62#, 8), to_unsigned(16#0E#, 8),
     to_unsigned(16#AA#, 8), to_unsigned(16#18#, 8), to_unsigned(16#BE#, 8), to_unsigned(16#1B#, 8),
     to_unsigned(16#FC#, 8), to_unsigned(16#56#, 8), to_unsigned(16#3E#, 8), to_unsigned(16#4B#, 8),
     to_unsigned(16#C6#, 8), to_unsigned(16#D2#, 8), to_unsigned(16#79#, 8), to_unsigned(16#20#, 8),
     to_unsigned(16#9A#, 8), to_unsigned(16#DB#, 8), to_unsigned(16#C0#, 8), to_unsigned(16#FE#, 8),
     to_unsigned(16#78#, 8), to_unsigned(16#CD#, 8), to_unsigned(16#5A#, 8), to_unsigned(16#F4#, 8),
     to_unsigned(16#1F#, 8), to_unsigned(16#DD#, 8), to_unsigned(16#A8#, 8), to_unsigned(16#33#, 8),
     to_unsigned(16#88#, 8), to_unsigned(16#07#, 8), to_unsigned(16#C7#, 8), to_unsigned(16#31#, 8),
     to_unsigned(16#B1#, 8), to_unsigned(16#12#, 8), to_unsigned(16#10#, 8), to_unsigned(16#59#, 8),
     to_unsigned(16#27#, 8), to_unsigned(16#80#, 8), to_unsigned(16#EC#, 8), to_unsigned(16#5F#, 8),
     to_unsigned(16#60#, 8), to_unsigned(16#51#, 8), to_unsigned(16#7F#, 8), to_unsigned(16#A9#, 8),
     to_unsigned(16#19#, 8), to_unsigned(16#B5#, 8), to_unsigned(16#4A#, 8), to_unsigned(16#0D#, 8),
     to_unsigned(16#2D#, 8), to_unsigned(16#E5#, 8), to_unsigned(16#7A#, 8), to_unsigned(16#9F#, 8),
     to_unsigned(16#93#, 8), to_unsigned(16#C9#, 8), to_unsigned(16#9C#, 8), to_unsigned(16#EF#, 8),
     to_unsigned(16#A0#, 8), to_unsigned(16#E0#, 8), to_unsigned(16#3B#, 8), to_unsigned(16#4D#, 8),
     to_unsigned(16#AE#, 8), to_unsigned(16#2A#, 8), to_unsigned(16#F5#, 8), to_unsigned(16#B0#, 8),
     to_unsigned(16#C8#, 8), to_unsigned(16#EB#, 8), to_unsigned(16#BB#, 8), to_unsigned(16#3C#, 8),
     to_unsigned(16#83#, 8), to_unsigned(16#53#, 8), to_unsigned(16#99#, 8), to_unsigned(16#61#, 8),
     to_unsigned(16#17#, 8), to_unsigned(16#2B#, 8), to_unsigned(16#04#, 8), to_unsigned(16#7E#, 8),
     to_unsigned(16#BA#, 8), to_unsigned(16#77#, 8), to_unsigned(16#D6#, 8), to_unsigned(16#26#, 8),
     to_unsigned(16#E1#, 8), to_unsigned(16#69#, 8), to_unsigned(16#14#, 8), to_unsigned(16#63#, 8),
     to_unsigned(16#55#, 8), to_unsigned(16#21#, 8), to_unsigned(16#0C#, 8), to_unsigned(16#7D#, 8));  -- ufix8 [256]
  CONSTANT nc_4                           : vector_of_unsigned8(0 TO 255) := 
    (to_unsigned(16#52#, 8), to_unsigned(16#09#, 8), to_unsigned(16#6A#, 8), to_unsigned(16#D5#, 8),
     to_unsigned(16#30#, 8), to_unsigned(16#36#, 8), to_unsigned(16#A5#, 8), to_unsigned(16#38#, 8),
     to_unsigned(16#BF#, 8), to_unsigned(16#40#, 8), to_unsigned(16#A3#, 8), to_unsigned(16#9E#, 8),
     to_unsigned(16#81#, 8), to_unsigned(16#F3#, 8), to_unsigned(16#D7#, 8), to_unsigned(16#FB#, 8),
     to_unsigned(16#7C#, 8), to_unsigned(16#E3#, 8), to_unsigned(16#39#, 8), to_unsigned(16#82#, 8),
     to_unsigned(16#9B#, 8), to_unsigned(16#2F#, 8), to_unsigned(16#FF#, 8), to_unsigned(16#87#, 8),
     to_unsigned(16#34#, 8), to_unsigned(16#8E#, 8), to_unsigned(16#43#, 8), to_unsigned(16#44#, 8),
     to_unsigned(16#C4#, 8), to_unsigned(16#DE#, 8), to_unsigned(16#E9#, 8), to_unsigned(16#CB#, 8),
     to_unsigned(16#54#, 8), to_unsigned(16#7B#, 8), to_unsigned(16#94#, 8), to_unsigned(16#32#, 8),
     to_unsigned(16#A6#, 8), to_unsigned(16#C2#, 8), to_unsigned(16#23#, 8), to_unsigned(16#3D#, 8),
     to_unsigned(16#EE#, 8), to_unsigned(16#4C#, 8), to_unsigned(16#95#, 8), to_unsigned(16#0B#, 8),
     to_unsigned(16#42#, 8), to_unsigned(16#FA#, 8), to_unsigned(16#C3#, 8), to_unsigned(16#4E#, 8),
     to_unsigned(16#08#, 8), to_unsigned(16#2E#, 8), to_unsigned(16#A1#, 8), to_unsigned(16#66#, 8),
     to_unsigned(16#28#, 8), to_unsigned(16#D9#, 8), to_unsigned(16#24#, 8), to_unsigned(16#B2#, 8),
     to_unsigned(16#76#, 8), to_unsigned(16#5B#, 8), to_unsigned(16#A2#, 8), to_unsigned(16#49#, 8),
     to_unsigned(16#6D#, 8), to_unsigned(16#8B#, 8), to_unsigned(16#D1#, 8), to_unsigned(16#25#, 8),
     to_unsigned(16#72#, 8), to_unsigned(16#F8#, 8), to_unsigned(16#F6#, 8), to_unsigned(16#64#, 8),
     to_unsigned(16#86#, 8), to_unsigned(16#68#, 8), to_unsigned(16#98#, 8), to_unsigned(16#16#, 8),
     to_unsigned(16#D4#, 8), to_unsigned(16#A4#, 8), to_unsigned(16#5C#, 8), to_unsigned(16#CC#, 8),
     to_unsigned(16#5D#, 8), to_unsigned(16#65#, 8), to_unsigned(16#B6#, 8), to_unsigned(16#92#, 8),
     to_unsigned(16#6C#, 8), to_unsigned(16#70#, 8), to_unsigned(16#48#, 8), to_unsigned(16#50#, 8),
     to_unsigned(16#FD#, 8), to_unsigned(16#ED#, 8), to_unsigned(16#B9#, 8), to_unsigned(16#DA#, 8),
     to_unsigned(16#5E#, 8), to_unsigned(16#15#, 8), to_unsigned(16#46#, 8), to_unsigned(16#57#, 8),
     to_unsigned(16#A7#, 8), to_unsigned(16#8D#, 8), to_unsigned(16#9D#, 8), to_unsigned(16#84#, 8),
     to_unsigned(16#90#, 8), to_unsigned(16#D8#, 8), to_unsigned(16#AB#, 8), to_unsigned(16#00#, 8),
     to_unsigned(16#8C#, 8), to_unsigned(16#BC#, 8), to_unsigned(16#D3#, 8), to_unsigned(16#0A#, 8),
     to_unsigned(16#F7#, 8), to_unsigned(16#E4#, 8), to_unsigned(16#58#, 8), to_unsigned(16#05#, 8),
     to_unsigned(16#B8#, 8), to_unsigned(16#B3#, 8), to_unsigned(16#45#, 8), to_unsigned(16#06#, 8),
     to_unsigned(16#D0#, 8), to_unsigned(16#2C#, 8), to_unsigned(16#1E#, 8), to_unsigned(16#8F#, 8),
     to_unsigned(16#CA#, 8), to_unsigned(16#3F#, 8), to_unsigned(16#0F#, 8), to_unsigned(16#02#, 8),
     to_unsigned(16#C1#, 8), to_unsigned(16#AF#, 8), to_unsigned(16#BD#, 8), to_unsigned(16#03#, 8),
     to_unsigned(16#01#, 8), to_unsigned(16#13#, 8), to_unsigned(16#8A#, 8), to_unsigned(16#6B#, 8),
     to_unsigned(16#3A#, 8), to_unsigned(16#91#, 8), to_unsigned(16#11#, 8), to_unsigned(16#41#, 8),
     to_unsigned(16#4F#, 8), to_unsigned(16#67#, 8), to_unsigned(16#DC#, 8), to_unsigned(16#EA#, 8),
     to_unsigned(16#97#, 8), to_unsigned(16#F2#, 8), to_unsigned(16#CF#, 8), to_unsigned(16#CE#, 8),
     to_unsigned(16#F0#, 8), to_unsigned(16#B4#, 8), to_unsigned(16#E6#, 8), to_unsigned(16#73#, 8),
     to_unsigned(16#96#, 8), to_unsigned(16#AC#, 8), to_unsigned(16#74#, 8), to_unsigned(16#22#, 8),
     to_unsigned(16#E7#, 8), to_unsigned(16#AD#, 8), to_unsigned(16#35#, 8), to_unsigned(16#85#, 8),
     to_unsigned(16#E2#, 8), to_unsigned(16#F9#, 8), to_unsigned(16#37#, 8), to_unsigned(16#E8#, 8),
     to_unsigned(16#1C#, 8), to_unsigned(16#75#, 8), to_unsigned(16#DF#, 8), to_unsigned(16#6E#, 8),
     to_unsigned(16#47#, 8), to_unsigned(16#F1#, 8), to_unsigned(16#1A#, 8), to_unsigned(16#71#, 8),
     to_unsigned(16#1D#, 8), to_unsigned(16#29#, 8), to_unsigned(16#C5#, 8), to_unsigned(16#89#, 8),
     to_unsigned(16#6F#, 8), to_unsigned(16#B7#, 8), to_unsigned(16#62#, 8), to_unsigned(16#0E#, 8),
     to_unsigned(16#AA#, 8), to_unsigned(16#18#, 8), to_unsigned(16#BE#, 8), to_unsigned(16#1B#, 8),
     to_unsigned(16#FC#, 8), to_unsigned(16#56#, 8), to_unsigned(16#3E#, 8), to_unsigned(16#4B#, 8),
     to_unsigned(16#C6#, 8), to_unsigned(16#D2#, 8), to_unsigned(16#79#, 8), to_unsigned(16#20#, 8),
     to_unsigned(16#9A#, 8), to_unsigned(16#DB#, 8), to_unsigned(16#C0#, 8), to_unsigned(16#FE#, 8),
     to_unsigned(16#78#, 8), to_unsigned(16#CD#, 8), to_unsigned(16#5A#, 8), to_unsigned(16#F4#, 8),
     to_unsigned(16#1F#, 8), to_unsigned(16#DD#, 8), to_unsigned(16#A8#, 8), to_unsigned(16#33#, 8),
     to_unsigned(16#88#, 8), to_unsigned(16#07#, 8), to_unsigned(16#C7#, 8), to_unsigned(16#31#, 8),
     to_unsigned(16#B1#, 8), to_unsigned(16#12#, 8), to_unsigned(16#10#, 8), to_unsigned(16#59#, 8),
     to_unsigned(16#27#, 8), to_unsigned(16#80#, 8), to_unsigned(16#EC#, 8), to_unsigned(16#5F#, 8),
     to_unsigned(16#60#, 8), to_unsigned(16#51#, 8), to_unsigned(16#7F#, 8), to_unsigned(16#A9#, 8),
     to_unsigned(16#19#, 8), to_unsigned(16#B5#, 8), to_unsigned(16#4A#, 8), to_unsigned(16#0D#, 8),
     to_unsigned(16#2D#, 8), to_unsigned(16#E5#, 8), to_unsigned(16#7A#, 8), to_unsigned(16#9F#, 8),
     to_unsigned(16#93#, 8), to_unsigned(16#C9#, 8), to_unsigned(16#9C#, 8), to_unsigned(16#EF#, 8),
     to_unsigned(16#A0#, 8), to_unsigned(16#E0#, 8), to_unsigned(16#3B#, 8), to_unsigned(16#4D#, 8),
     to_unsigned(16#AE#, 8), to_unsigned(16#2A#, 8), to_unsigned(16#F5#, 8), to_unsigned(16#B0#, 8),
     to_unsigned(16#C8#, 8), to_unsigned(16#EB#, 8), to_unsigned(16#BB#, 8), to_unsigned(16#3C#, 8),
     to_unsigned(16#83#, 8), to_unsigned(16#53#, 8), to_unsigned(16#99#, 8), to_unsigned(16#61#, 8),
     to_unsigned(16#17#, 8), to_unsigned(16#2B#, 8), to_unsigned(16#04#, 8), to_unsigned(16#7E#, 8),
     to_unsigned(16#BA#, 8), to_unsigned(16#77#, 8), to_unsigned(16#D6#, 8), to_unsigned(16#26#, 8),
     to_unsigned(16#E1#, 8), to_unsigned(16#69#, 8), to_unsigned(16#14#, 8), to_unsigned(16#63#, 8),
     to_unsigned(16#55#, 8), to_unsigned(16#21#, 8), to_unsigned(16#0C#, 8), to_unsigned(16#7D#, 8));  -- ufix8 [256]
END mlhdlc_aesd_fixpt_pkg;




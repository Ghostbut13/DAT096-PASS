-------------------------------------------------------------------------------
-- Title      : Wrapper ---- Config-i2c (ACFC-I2C)
-- Project    : 
-------------------------------------------------------------------------------
-- File       : Wrapper-ACFC_i2c.vhdl
-- Author     : Weihan Gao -- weihanga@chalmers.se
-- Company    : 
-- Created    : 2023-02-08
-- Last update: 2023-02-11
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: 
-------------------------------------------------------------------------------
-- Copyright (c) 2023 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2023-02-08  1.0      ASUS	Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Wrapper_ACFC_i2c is

  GENERIC(WORD_LENGHT: NATURAL RANGE 1 TO 128 := 16) ;
  port (
    -- finish config
    finish_config_input : in std_logic;
    -- CONfig THE MODE
    I2S_mode    : in  std_logic;
    master_mode : in  std_logic;
    GPIO_MCLK   : in  std_logic;
    FS_48k_256_BCLK  : in  std_logic;
    MCLK_root  : in std_logic;

    -- MCLK(GPIO)-generated by PLL and SHDNZ
    SHDNZ     : out    std_logic;
    MCLK      : out    std_logic;

    -- clk and rstn
    clk       : in    std_logic;
    rstn      : in    std_logic;
    -- control ready
    SW_vdd_ok : in    std_logic;
    SHDNZ_ready : in    std_logic;
    
    -- FSYNC and BCLK 
    FSYNC     : in   std_logic;
    BCLK      : in   std_logic;
    
    -- i2c communication
    SDA       : inout std_logic;
    SCL       : out   std_logic;
    
	--i2s communication
	DIN : in std_logic;
	start_I2S : in std_logic; 
	L1_out : out std_logic_vector (WORD_LENGHT-1 downto 0)
--	L2_out : out std_logic_vector (WORD_LENGHT-1 downto 0);
--	R1_out : out std_logic_vector (WORD_LENGHT-1 downto 0);
--	R2_out : out std_logic_vector (WORD_LENGHT-1 downto 0)
    );

end entity Wrapper_ACFC_i2c;


architecture arch_Wrapper_ACFC_i2c of Wrapper_ACFC_i2c is
  -- component
  component ADC_Configuration_Flow_Controller is
    -- generic(
    --   -- MODE reg addr
    --   constant const_addr_sleep_reg         : std_logic_vector(7 downto 0) := x"02";
    --   constant const_addr_interrupt_reg     : std_logic_vector(7 downto 0) := x"28";
    --   constant const_addr_c1_reg            : std_logic_vector(7 downto 0) := x"3c";
    --   constant const_addr_c2_reg            : std_logic_vector(7 downto 0) := x"41";
    --   constant const_addr_c3_reg            : std_logic_vector(7 downto 0) := x"46";
    --   constant const_addr_c4_reg            : std_logic_vector(7 downto 0) := x"4b";
    --   constant const_addr_input_channel_reg : std_logic_vector(7 downto 0) := x"73";
    --   constant const_addr_8_reg             : std_logic_vector(7 downto 0) := x"74";
    --   constant const_addr_powerup_reg       : std_logic_vector(7 downto 0) := x"75";
    --   constant const_addr_10_reg            : std_logic_vector(7 downto 0) := x"64"
    --   );
    port (
      finish_config_input : in std_logic;
      I2S_mode    : in  std_logic;
      master_mode : in  std_logic;
      GPIO_MCLK   : in  std_logic;
      FS_48k_256_BCLK  : in  std_logic;
      MCLK_root  : in std_logic;
      
      rstn         : in  std_logic;
      clk          : in  std_logic;
      done         : in  std_logic;
      start        : out std_logic;
      config_value : out std_logic_vector(7 downto 0);
      config_addr  : out std_logic_vector(7 downto 0);
      SHDNZ        : out std_logic;
      SHDNZ_ready  : in  std_logic;
      SW_vdd_ok    : in  std_logic
      );
  end component ADC_Configuration_Flow_Controller;
  
  component I2C_Interface is
    port (
      clk  : in std_logic;
      rstn : in std_logic;
      -- signals between i2c and ACFC
      start : in std_logic;
      done : out std_logic;
      config_addr : in  std_logic_vector(7 downto 0);
      config_value : in  std_logic_vector(7 downto 0);
      -- i2c communication
      SDA : inout std_logic;
      SCL : out std_logic
      );
  end component I2C_Interface;

---------------------
  component PLL_12M is
 port (
    clk_out1_0 : out STD_LOGIC;
    reset : in STD_LOGIC;
    sys_clock : in STD_LOGIC
  );
  end component PLL_12M;

  ------------------------------------------------------------
  -- signal between i2c and ACFC
  signal done : std_logic;
  signal start : std_logic;
  signal config_value : std_logic_vector(7 downto 0);
  signal config_addr  : std_logic_vector(7 downto 0);
  -- out signal for FSYNC and BCLK
  signal out_FSYNC : std_logic;
  signal out_BCLK : std_logic;

  signal out_n_clk : std_logic;
  signal out_p_clk : std_logic;
  
	signal L1_signal :  std_logic_vector (WORD_LENGHT-1 downto 0);
	signal	L2_signal :  std_logic_vector (WORD_LENGHT-1 downto 0);
	signal	R1_signal :  std_logic_vector (WORD_LENGHT-1 downto 0);
	signal	R2_signal :  std_logic_vector (WORD_LENGHT-1 downto 0);

  

component I2S IS
 GENERIC(WORD_LENGHT: NATURAL RANGE 1 TO 128) ;
 PORT  (
		bclk:IN STD_LOGIC ;
		start:IN STD_LOGIC ;
		reset:IN STD_LOGIC ;
		fsync:IN STD_LOGIC ;
		DIN : IN STD_LOGIC;
		LC_1_out : out std_logic_vector (WORD_LENGHT-1 downto 0)
--		LC_2_out : out std_logic_vector (WORD_LENGHT-1 downto 0);
--		RC_1_out : out std_logic_vector (WORD_LENGHT-1 downto 0);
--		RC_2_out : out std_logic_vector (WORD_LENGHT-1 downto 0);
--		SDOUT : OUT std_logic
		);
END component I2S;



  
    
begin  -- architecture arch_Wrapper_ACFC_i2c
  
  --FSYNC <=  out_FSYNC;
  --BCLK <=  out_BCLK;

  out_p_clk <= not(out_n_clk);
  out_n_clk <= clk;
  
  ------------------------------------------------------------
  -- INSTANCE
  inst_ACFC: component ADC_Configuration_Flow_Controller
    port map (
      finish_config_input => finish_config_input,
      I2S_mode     => I2S_mode,
      master_mode  => master_mode,
      GPIO_MCLK    => GPIO_MCLK  ,
      FS_48k_256_BCLK   => FS_48k_256_BCLK,
      MCLK_root  => MCLK_root,

      rstn         => rstn,
      clk          => clk,
      done         => done,
      start        => start,
      config_value => config_value,
      config_addr  => config_addr,
      SHDNZ        => SHDNZ,
      SHDNZ_ready  => SHDNZ_ready,
      SW_vdd_ok    => SW_vdd_ok);
  inst_i2c: component I2C_Interface
    port map (
      clk   => clk,
      rstn  => rstn,
      config_addr => config_addr,
      config_value => config_value,
      start => start,
      done  => done,
      SDA   => SDA,
      SCL   => SCL );
  inst_i2S: component I2S
  
    generic map (WORD_LENGHT=>WORD_LENGHT)
    port map (
    bclk =>BCLK,
	start =>start_I2S,
	reset =>rstn,
	fsync =>FSYNC,
	DIN =>DIN,
	LC_1_out => L1_signal);
		
--	LC_2_out =>L2_signal,
--	RC_1_out =>R1_signal,
--	RC_2_out =>  R2_signal);
      
  ------------------------------------------------------------
  ----GENERATE the FSYNC and BCLK by PLL
clk_wiz_0: component PLL_12M
     port map (
     sys_clock => clk,
      clk_out1_0 => MCLK,
      reset => rstn
    );
  ------------------------------------------------------------
  
  
end architecture arch_Wrapper_ACFC_i2c;
